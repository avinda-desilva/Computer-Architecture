//implement your 32-bit ALU
module alu32(out, overflow, zero, negative, A, B, control);
    output [31:0] out;
    output        overflow, zero, negative;
    input  [31:0] A, B;
    input   [2:0] control;
    wire [31:0] cin_in;
    wire [30:0] chain;
    wire cout;

    alu1 a1(out[0], cin_in[0], A[0], B[0], control[0], control);
    alu1 a2(out[1], cin_in[1], A[1], B[1], cin_in[0], control);
    alu1 a3(out[2], cin_in[2], A[2], B[2], cin_in[1], control);
    alu1 a4(out[3], cin_in[3], A[3], B[3], cin_in[2], control);
    alu1 a5(out[4], cin_in[4], A[4], B[4], cin_in[3], control);
    alu1 a6(out[5], cin_in[5], A[5], B[5], cin_in[4], control);
    alu1 a7(out[6], cin_in[6], A[6], B[6], cin_in[5], control);
    alu1 a8(out[7], cin_in[7], A[7], B[7], cin_in[6], control);
    alu1 a9(out[8], cin_in[8], A[8], B[8], cin_in[7], control);
    alu1 a10(out[9], cin_in[9], A[9], B[9], cin_in[8], control);
    alu1 a11(out[10], cin_in[10], A[10], B[10], cin_in[9], control);
    alu1 a12(out[11], cin_in[11], A[11], B[11], cin_in[10], control);
    alu1 a13(out[12], cin_in[12], A[12], B[12], cin_in[11], control);
    alu1 a14(out[13], cin_in[13], A[13], B[13], cin_in[12], control);
    alu1 a15(out[14], cin_in[14], A[14], B[14], cin_in[13], control);
    alu1 a16(out[15], cin_in[15], A[15], B[15], cin_in[14], control);
    alu1 a17(out[16], cin_in[16], A[16], B[16], cin_in[15], control);
    alu1 a18(out[17], cin_in[17], A[17], B[17], cin_in[16], control);
    alu1 a19(out[18], cin_in[18], A[18], B[18], cin_in[17], control);
    alu1 a20(out[19], cin_in[19], A[19], B[19], cin_in[18], control);
    alu1 a21(out[20], cin_in[20], A[20], B[20], cin_in[19], control);
    alu1 a22(out[21], cin_in[21], A[21], B[21], cin_in[20], control);
    alu1 a23(out[22], cin_in[22], A[22], B[22], cin_in[21], control);
    alu1 a24(out[23], cin_in[23], A[23], B[23], cin_in[22], control);
    alu1 a25(out[24], cin_in[24], A[24], B[24], cin_in[23], control);
    alu1 a26(out[25], cin_in[25], A[25], B[25], cin_in[24], control);
    alu1 a27(out[26], cin_in[26], A[26], B[26], cin_in[25], control);
    alu1 a28(out[27], cin_in[27], A[27], B[27], cin_in[26], control);
    alu1 a29(out[28], cin_in[28], A[28], B[28], cin_in[27], control);
    alu1 a30(out[29], cin_in[29], A[29], B[29], cin_in[28], control);
    alu1 a31(out[30], cin_in[30], A[30], B[30], cin_in[29], control);
    alu1 a32(out[31], cin_in[31], A[31], B[31], cin_in[30], control);

    assign negative = out[31];
    or o1(chain[0], out[1], out[0]);
    or o2(chain[1], out[2], chain[0]);
    or o3(chain[2], out[3], chain[1]);
    or o4(chain[3], out[4], chain[2]);
    or o5(chain[4], out[5], chain[3]);
    or o6(chain[5], out[6], chain[4]);
    or o7(chain[6], out[7], chain[5]);
    or o8(chain[7], out[8], chain[6]);
    or o9(chain[8], out[9], chain[7]);
    or o10(chain[9], out[10], chain[8]);
    or o11(chain[10], out[11], chain[9]);
    or o12(chain[11], out[12], chain[10]);
    or o13(chain[12], out[13], chain[11]);
    or o14(chain[13], out[14], chain[12]);
    or o15(chain[14], out[15], chain[13]);
    or o16(chain[15], out[16], chain[14]);
    or o17(chain[16], out[17], chain[15]);
    or o18(chain[17], out[18], chain[16]);
    or o19(chain[18], out[19], chain[17]);
    or o20(chain[19], out[20], chain[18]);
    or o21(chain[20], out[21], chain[19]);
    or o22(chain[21], out[22], chain[20]);
    or o23(chain[22], out[23], chain[21]);
    or o24(chain[23], out[24], chain[22]);
    or o25(chain[24], out[25], chain[23]);
    or o26(chain[25], out[26], chain[24]);
    or o27(chain[26], out[27], chain[25]);
    or o28(chain[27], out[28], chain[26]);
    or o29(chain[28], out[29], chain[27]);
    or o30(chain[29], out[30], chain[28]);
    or o31(chain[30], out[31], chain[29]);
    not n1(zero, chain[30]);
    xor x1(overflow, cin_in[31], cin_in[30]);

endmodule // alu32
